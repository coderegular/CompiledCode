AND(a,b,c)
OR(x,y,z)
NOT(b,y)
NAND(c,d,b)
NOR(z,t,b)
XOR(t,a,x)
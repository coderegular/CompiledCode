AND(e,a,b)
OR(h,c,d)
OR(k,e,h)
AND(l,e,h)
OR(t,c,d)
NAND(p,k,l)
